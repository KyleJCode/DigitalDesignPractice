module RRPolicy();
// Replaces random block in memory.



endmodule
module LFUPolicy();
// Replaces the least frequently used block in memory.



endmodule
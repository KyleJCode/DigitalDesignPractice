module LRUPolicy();
// Replaces the least recently used block in memory.


endmodule
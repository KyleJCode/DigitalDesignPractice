module LRUPolicy();
// Replaces the least recently used block in memory. Essentially a FIFO.


endmodule
module DataLogger(rst, clk, policy_sel, log_en,);



endmodule
module SizePolicy();
// Replaces largest sized block in memory.



endmodule